// riscxv_top_tb.sv
module riscxv_top_tb;

    // Input and output ports can be left empty for now

    initial begin
        $display("Testbench for riscxv started.");
        // Add simulation initialization here
    end

endmodule
