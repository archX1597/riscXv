// riscxv_pkg.sv
package riscxv_pkg;

    // Define common types, parameters, and constants here

endpackage
